`timescale 1ns / 1ps

module soc_top
  (
    input wire [31:0]  saxi_araddr,
    input wire [1:0]   saxi_arburst,
    input wire [3:0]   saxi_arcache,
    input wire [3:0]   saxi_arid,
    input wire [7:0]   saxi_arlen,
    input wire         saxi_arlock,
    input wire [2:0]   saxi_arprot,
    input wire [3:0]   saxi_arqos,
    input wire [3:0]   saxi_arregion,
    input wire [2:0]   saxi_arsize,
    output wire        saxi_arready,
    input wire         saxi_arvalid,
    input wire [31:0]  saxi_awaddr,
    input wire [1:0]   saxi_awburst,
    input wire [3:0]   saxi_awcache,
    input wire [3:0]   saxi_awid,
    input wire [7:0]   saxi_awlen,
    input wire         saxi_awlock,
    input wire [2:0]   saxi_awprot,
    input wire [3:0]   saxi_awqos,
    input wire [3:0]   saxi_awregion,
    input wire [2:0]   saxi_awsize,
    output wire        saxi_awready,
    input wire         saxi_awvalid,
    output wire [3:0]  saxi_bid,
    output wire [1:0]  saxi_bresp,
    input wire         saxi_bready,
    output wire        saxi_bvalid,
    output wire [63:0] saxi_rdata,
    output wire [3:0]  saxi_rid,
    output wire        saxi_rlast,
    output wire [1:0]  saxi_rresp,
    input wire         saxi_rready,
    output wire        saxi_rvalid,
    input wire [63:0]  saxi_wdata,
    input wire         saxi_wlast,
    input wire [7:0]   saxi_wstrb,
    output wire        saxi_wready,
    input wire         saxi_wvalid,
    input wire [31:0]  saxil_araddr,
    input wire [2:0]   saxil_arprot,
    output wire        saxil_arready,
    input wire         saxil_arvalid,
    input wire [31:0]  saxil_awaddr,
    input wire [2:0]   saxil_awprot,
    output wire        saxil_awready,
    input wire         saxil_awvalid,
    input wire         saxil_bready,
    output wire [1:0]  saxil_bresp,
    output wire        saxil_bvalid,
    output wire [31:0] saxil_rdata,
    input wire         saxil_rready,
    output wire [1:0]  saxil_rresp,
    output wire        saxil_rvalid,
    input wire [31:0]  saxil_wdata,
    output wire        saxil_wready,
    input wire [3:0]   saxil_wstrb,
    input wire         saxil_wvalid,
    output wire [29:0] maxi_araddr,
    output wire [1:0]  maxi_arburst,
    output wire [3:0]  maxi_arcache,
    output wire [5:0]  maxi_arid,
    output wire [7:0]  maxi_arlen,
    output wire        maxi_arlock,
    output wire [2:0]  maxi_arprot,
    output wire [3:0]  maxi_arqos,
    output wire [3:0]  maxi_arregion,
    output wire [2:0]  maxi_arsize,
    input wire         maxi_arready,
    output wire        maxi_arvalid,
    output wire [29:0] maxi_awaddr,
    output wire [1:0]  maxi_awburst,
    output wire [3:0]  maxi_awcache,
    output wire [5:0]  maxi_awid,
    output wire [7:0]  maxi_awlen,
    output wire        maxi_awlock,
    output wire [2:0]  maxi_awprot,
    output wire [3:0]  maxi_awqos,
    output wire [3:0]  maxi_awregion,
    output wire [2:0]  maxi_awsize,
    input wire         maxi_awready,
    output wire        maxi_awvalid,
    input wire [5:0]   maxi_bid,
    input wire [1:0]   maxi_bresp,
    output wire        maxi_bready,
    input wire         maxi_bvalid,
    input wire [63:0]  maxi_rdata,
    input wire [5:0]   maxi_rid,
    input wire         maxi_rlast,
    input wire [1:0]   maxi_rresp,
    output wire        maxi_rready,
    input wire         maxi_rvalid,
    output wire [63:0] maxi_wdata,
    output wire        maxi_wlast,
    output wire [7:0]  maxi_wstrb,
    input wire         maxi_wready,
    output wire        maxi_wvalid,
    input wire         uart_rx,
    output wire        uart_tx,
    output wire        sdio_ck,
    inout wire         sdio_cmd,
    inout wire [3:0]   sdio_data,
    input              clk,
    input              aresetn
   );

   wire                         jtag_tck;
   wire                         jtag_tdi;
   wire                         jtag_tms;
   wire                         jtag_tdo;

   JTAGTUNNEL jtagtunnel
     (
      .jtag_tck(jtag_tck),
      .jtag_tdi(jtag_tdi),
      .jtag_tms(jtag_tms),
      .jtag_tdo(jtag_tdo),
      .jtag_tdo_en(1'b1)
      );

   wire                         sdio_cmd_i;
   wire                         sdio_cmd_o;
   wire                         sdio_cmt_t;

   wire [3:0]                   sdio_data_i;
   wire [3:0]                   sdio_data_o;
   wire [3:0]                   sdio_data_t;

   IOBUF #(.IOSTANDARD("LVCMOS33"))
   IOBUF_cmd(
             .O(sdio_cmd_i),
             .IO(sdio_cmd),
             .I(sdio_cmd_o),
             .T(sdio_cmd_t)
             );

   genvar                       i;
   generate
      for (i = 0; i < 4; i = i+1) begin
         IOBUF #(.IOSTANDARD("LVCMOS33"))
         IOBUF_data
           (
            .O(sdio_data_i[i]),
            .IO(sdio_data[i]),
            .I(sdio_data_o[i]),
            .T(sdio_data_t[i])
            );
      end
   endgenerate

   soc_wrapper soc_wrapper
     (
      .axi_master__ar__bits__addr(saxi_araddr),
      .axi_master__ar__bits__burst(saxi_arburst),
      .axi_master__ar__bits__cache(saxi_arcache),
      .axi_master__ar__bits__id(saxi_arid),
      .axi_master__ar__bits__len(saxi_arlen),
      .axi_master__ar__bits__lock(saxi_arlock),
      .axi_master__ar__bits__prot(saxi_arprot),
      .axi_master__ar__bits__qos(saxi_arqos),
      .axi_master__ar__bits__region(saxi_arregion),
      .axi_master__ar__bits__size(saxi_arsize),
      .axi_master__ar__ready(saxi_arready),
      .axi_master__ar__valid(saxi_arvalid),
      .axi_master__aw__bits__addr(saxi_awaddr),
      .axi_master__aw__bits__burst(saxi_awburst),
      .axi_master__aw__bits__cache(saxi_awcache),
      .axi_master__aw__bits__id(saxi_awid),
      .axi_master__aw__bits__len(saxi_awlen),
      .axi_master__aw__bits__lock(saxi_awlock),
      .axi_master__aw__bits__prot(saxi_awprot),
      .axi_master__aw__bits__qos(saxi_awqos),
      .axi_master__aw__bits__region(saxi_awregion),
      .axi_master__aw__bits__size(saxi_awsize),
      .axi_master__aw__ready(saxi_awready),
      .axi_master__aw__valid(saxi_awvalid),
      .axi_master__b__bits__id(saxi_bid),
      .axi_master__b__bits__resp(saxi_bresp),
      .axi_master__b__ready(saxi_bready),
      .axi_master__b__valid(saxi_bvalid),
      .axi_master__r__bits__data(saxi_rdata),
      .axi_master__r__bits__id(saxi_rid),
      .axi_master__r__bits__last(saxi_rlast),
      .axi_master__r__bits__resp(saxi_rresp),
      .axi_master__r__ready(saxi_rready),
      .axi_master__r__valid(saxi_rvalid),
      .axi_master__w__bits__data(saxi_wdata),
      .axi_master__w__bits__last(saxi_wlast),
      .axi_master__w__bits__strb(saxi_wstrb),
      .axi_master__w__ready(saxi_wready),
      .axi_master__w__valid(saxi_wvalid),
      .axil_master__ar__addr(saxil_araddr),
      .axil_master__ar__prot(saxil_arprot),
      .axil_master__ar__ready(saxil_arready),
      .axil_master__ar__valid(saxil_arvalid),
      .axil_master__aw__addr(saxil_awaddr),
      .axil_master__aw__prot(saxil_awprot),
      .axil_master__aw__ready(saxil_awready),
      .axil_master__aw__valid(saxil_awvalid),
      .axil_master__b__ready(saxil_bready),
      .axil_master__b__resp(saxil_bresp),
      .axil_master__b__valid(saxil_bvalid),
      .axil_master__r__data(saxil_rdata),
      .axil_master__r__ready(saxil_rready),
      .axil_master__r__resp(saxil_rresp),
      .axil_master__r__valid(saxil_rvalid),
      .axil_master__w__data(saxil_wdata),
      .axil_master__w__ready(saxil_wready),
      .axil_master__w__strb(saxil_wstrb),
      .axil_master__w__valid(saxil_wvalid),
      .ram_bus__ar__bits__addr(maxi_araddr),
      .ram_bus__ar__bits__burst(maxi_arburst),
      .ram_bus__ar__bits__cache(maxi_arcache),
      .ram_bus__ar__bits__id(maxi_arid),
      .ram_bus__ar__bits__len(maxi_arlen),
      .ram_bus__ar__bits__lock(maxi_arlock),
      .ram_bus__ar__bits__prot(maxi_arprot),
      .ram_bus__ar__bits__qos(maxi_arqos),
      .ram_bus__ar__bits__region(maxi_arregion),
      .ram_bus__ar__bits__size(maxi_arsize),
      .ram_bus__ar__ready(maxi_arready),
      .ram_bus__ar__valid(maxi_arvalid),
      .ram_bus__aw__bits__addr(maxi_awaddr),
      .ram_bus__aw__bits__burst(maxi_awburst),
      .ram_bus__aw__bits__cache(maxi_awcache),
      .ram_bus__aw__bits__id(maxi_awid),
      .ram_bus__aw__bits__len(maxi_awlen),
      .ram_bus__aw__bits__lock(maxi_awlock),
      .ram_bus__aw__bits__prot(maxi_awprot),
      .ram_bus__aw__bits__qos(maxi_awqos),
      .ram_bus__aw__bits__region(maxi_awregion),
      .ram_bus__aw__bits__size(maxi_awsize),
      .ram_bus__aw__ready(maxi_awready),
      .ram_bus__aw__valid(maxi_awvalid),
      .ram_bus__b__bits__id(maxi_bid),
      .ram_bus__b__bits__resp(maxi_bresp),
      .ram_bus__b__ready(maxi_bready),
      .ram_bus__b__valid(maxi_bvalid),
      .ram_bus__r__bits__data(maxi_rdata),
      .ram_bus__r__bits__id(maxi_rid),
      .ram_bus__r__bits__last(maxi_rlast),
      .ram_bus__r__bits__resp(maxi_rresp),
      .ram_bus__r__ready(maxi_rready),
      .ram_bus__r__valid(maxi_rvalid),
      .ram_bus__w__bits__data(maxi_wdata),
      .ram_bus__w__bits__last(maxi_wlast),
      .ram_bus__w__bits__strb(maxi_wstrb),
      .ram_bus__w__ready(maxi_wready),
      .ram_bus__w__valid(maxi_wvalid),
      .tck(jtag_tck),
      .tdi(jtag_tdi),
      .tms(jtag_tms),
      .tdo(jtag_tdo),
      .rx(uart_rx),
      .tx(uart_tx),
      .sdio_clk(sdio_ck),
      .sdio_cmd_i(sdio_cmd_i),
      .sdio_cmd_o(sdio_cmd_o),
      .sdio_cmd_t(sdio_cmd_t),
      .sdio_data_i(sdio_data_i),
      .sdio_data_o(sdio_data_o),
      .sdio_data_t(sdio_data_t),
      .clk(clk),
      .rst(~aresetn)
      );

endmodule
